module dcache (
    input
